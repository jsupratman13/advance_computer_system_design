library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.led_matrix.all;

entity ART is
    port(
        FLAG      : in integer;
        GRID      : out std_matrix);
end ART;

architecture RTL of ART is
    signal NO_ART   : std_matrix := ((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

    signal ART0   : std_matrix :=   ((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3),
                                     (3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3),
                                     (3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3),
                                     (3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3),
                                     (3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3),
                                     (3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3),
                                     (3,3,3,3,3,3,3,3,3,3,3,3,3,3,3,3),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

    signal ART1     : std_matrix := ((0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,1,1,1,1,0,0,0,0,0,0),
                                     (0,0,0,0,0,1,1,0,1,1,0,0,0,0,0,0),
                                     (0,0,0,0,0,1,0,0,1,1,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0),
                                     (0,0,0,1,1,1,1,1,1,1,1,1,1,1,0,0),
                                     (0,0,0,1,1,1,1,1,1,1,1,1,1,1,0,0));

    signal ART2     : std_matrix := ((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
                                     (1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
                                     (1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

    signal ART3   : std_matrix :=   ((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
                                     (2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
                                     (2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
                                     (2,2,2,2,2,2,2,2,2,2,2,2,2,2,2,2),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                     (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

    begin
        process(FLAG) begin
            case FLAG is
                when 0 => GRID <= ART0;
                when 1 => GRID <= ART1;
                when 2 => GRID <= ART2;
                when 3 => GRID <= ART3;
                when others => GRID <= NO_ART;
				end case;
        end process;

end RTL;
        
