library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.led_matrix.all;

entity ART is
    port(
        FLAG      : in integer;
        GRID      : out std_matrix);
end ART;

architecture RTL of ART is
    constant NO_ART   : std_matrix := ((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

    constant ART0     : std_matrix := ((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0),
                                       (0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0),
                                       (0,0,0,0,0,0,1,0,0,0,1,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,1,0,1,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

    constant ART1     : std_matrix := ((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,2,2,2,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,2,0,0,0,2,0,0,0,0),
                                       (0,0,0,0,0,0,2,0,0,0,0,0,2,0,0,0),
                                       (0,0,0,0,0,0,2,0,0,0,0,0,2,0,0,0),
                                       (0,0,0,0,0,0,2,0,0,0,0,0,2,0,0,0),
                                       (0,0,0,0,0,0,0,2,0,0,0,0,2,0,0,0),
                                       (0,0,0,0,0,0,0,0,2,0,0,2,2,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,2,2,0,2,0,0,0),
                                       (0,0,0,0,0,0,0,0,2,0,0,0,2,0,0,0),
                                       (0,0,0,0,0,0,0,2,0,0,0,0,2,0,0,0),
                                       (0,0,0,0,0,0,2,0,0,0,0,0,2,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

    constant ART2     : std_matrix := ((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,2,2,2,2,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,2,2,2,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

    constant ART3     : std_matrix := ((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,2,2,2,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,2,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,2,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,2,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,2,2,2,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));


    constant ART4     : std_matrix := ((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,2,2,2,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,2,2,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,2,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,2,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,2,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,2,2,2,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

    constant ART5     : std_matrix := ((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,2,2,2,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,2,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,2,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,2,2,2,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,2,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,2,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,2,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,2,0,0,0,2,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

    constant ART6     : std_matrix := ((0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,1,1,0,0,0,0,1,1,0,0,0,0),
                                       (0,0,0,1,0,0,2,0,0,2,0,0,1,0,0,0),
                                       (0,0,1,0,0,0,2,0,0,2,0,0,0,1,0,0),
                                       (0,0,1,0,0,0,0,2,2,0,0,0,0,1,0,0),
                                       (0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0),
                                       (0,0,0,0,1,2,0,0,0,0,2,1,0,0,0,0),
                                       (0,0,0,0,0,1,0,0,0,0,1,0,0,0,0,0),
                                       (0,0,0,0,0,1,0,0,0,0,1,0,0,0,0,0),
                                       (0,0,0,0,0,0,1,0,0,1,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
                                       (0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0));

    begin
        process(FLAG) begin
            case FLAG is
                when 0 => GRID <= ART0;
                when 1 => GRID <= ART1;
                when 2 => GRID <= ART2;
                when 3 => GRID <= ART3;
                when 4 => GRID <= ART4;
                when 5 => GRID <= ART5;
                when 6 => GRID <= ART6;
                when others => GRID <= NO_ART;
				end case;
        end process;

end RTL;
        
